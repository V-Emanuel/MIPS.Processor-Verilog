module Module_AND (ent1, ent2, saida);

	input ent1, ent2;
	output saida;
	assign saida = ent1 & ent2;
	
endmodule
